library verilog;
use verilog.vl_types.all;
entity ControleTemp_vlg_vec_tst is
end ControleTemp_vlg_vec_tst;
